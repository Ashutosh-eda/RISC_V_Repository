// ============================================================================
// Leading Zero Counter (LZC)
// Uses priority encoder to count leading zeros in a 48-bit value
// Critical for normalization shift amount calculation
// ============================================================================

module fpu_lzc (
    input  wire [47:0] data_in,
    output reg  [5:0]  count       // 0-48 leading zeros
);

    // Priority encoder - find first '1' bit from MSB
    always @(*) begin
        casez (data_in)
            48'b1???????????????????????????????????????????????: count = 6'd0;
            48'b01??????????????????????????????????????????????: count = 6'd1;
            48'b001?????????????????????????????????????????????: count = 6'd2;
            48'b0001????????????????????????????????????????????: count = 6'd3;
            48'b00001???????????????????????????????????????????: count = 6'd4;
            48'b000001??????????????????????????????????????????: count = 6'd5;
            48'b0000001?????????????????????????????????????????: count = 6'd6;
            48'b00000001????????????????????????????????????????: count = 6'd7;
            48'b000000001???????????????????????????????????????: count = 6'd8;
            48'b0000000001??????????????????????????????????????: count = 6'd9;
            48'b00000000001?????????????????????????????????????: count = 6'd10;
            48'b000000000001????????????????????????????????????: count = 6'd11;
            48'b0000000000001???????????????????????????????????: count = 6'd12;
            48'b00000000000001??????????????????????????????????: count = 6'd13;
            48'b000000000000001?????????????????????????????????: count = 6'd14;
            48'b0000000000000001????????????????????????????????: count = 6'd15;
            48'b00000000000000001???????????????????????????????: count = 6'd16;
            48'b000000000000000001??????????????????????????????: count = 6'd17;
            48'b0000000000000000001?????????????????????????????: count = 6'd18;
            48'b00000000000000000001????????????????????????????: count = 6'd19;
            48'b000000000000000000001???????????????????????????: count = 6'd20;
            48'b0000000000000000000001??????????????????????????: count = 6'd21;
            48'b00000000000000000000001?????????????????????????: count = 6'd22;
            48'b000000000000000000000001????????????????????????: count = 6'd23;
            48'b0000000000000000000000001???????????????????????: count = 6'd24;
            48'b00000000000000000000000001??????????????????????: count = 6'd25;
            48'b000000000000000000000000001?????????????????????: count = 6'd26;
            48'b0000000000000000000000000001????????????????????: count = 6'd27;
            48'b00000000000000000000000000001???????????????????: count = 6'd28;
            48'b000000000000000000000000000001??????????????????: count = 6'd29;
            48'b0000000000000000000000000000001?????????????????: count = 6'd30;
            48'b00000000000000000000000000000001????????????????: count = 6'd31;
            48'b000000000000000000000000000000001???????????????: count = 6'd32;
            48'b0000000000000000000000000000000001??????????????: count = 6'd33;
            48'b00000000000000000000000000000000001?????????????: count = 6'd34;
            48'b000000000000000000000000000000000001????????????: count = 6'd35;
            48'b0000000000000000000000000000000000001???????????: count = 6'd36;
            48'b00000000000000000000000000000000000001??????????: count = 6'd37;
            48'b000000000000000000000000000000000000001?????????: count = 6'd38;
            48'b0000000000000000000000000000000000000001????????: count = 6'd39;
            48'b00000000000000000000000000000000000000001???????: count = 6'd40;
            48'b000000000000000000000000000000000000000001??????: count = 6'd41;
            48'b0000000000000000000000000000000000000000001?????: count = 6'd42;
            48'b00000000000000000000000000000000000000000001????: count = 6'd43;
            48'b000000000000000000000000000000000000000000001???: count = 6'd44;
            48'b0000000000000000000000000000000000000000000001??: count = 6'd45;
            48'b00000000000000000000000000000000000000000000001?: count = 6'd46;
            48'b000000000000000000000000000000000000000000000001: count = 6'd47;
            48'b000000000000000000000000000000000000000000000000: count = 6'd48;  // All zeros
            default: count = 6'd0;
        endcase
    end

endmodule
